`timescale 1ns / 1ps
module InstMem(Address, Instruction);
    input wire [31:0] Address;
	output reg [31:0] Instruction;

	parameter MEM_SIZE = 512;
	reg [31:0] data [MEM_SIZE - 1:0];	

    //assign Instruction = data[Address[10:2]];
    
    always @(*) begin
        case(Address[10:2])
        9'd0	:	 Instruction <= 32'h20040006	;
        9'd1    :    Instruction <= 32'hac040000    ;
        9'd2    :    Instruction <= 32'h20050004    ;
        9'd3    :    Instruction <= 32'h20060320    ;
        9'd4    :    Instruction <= 32'h20070348    ;
        9'd5    :    Instruction <= 32'h20a90000    ;
        9'd6    :    Instruction <= 32'h24080000    ;
        9'd7    :    Instruction <= 32'had280000    ;
        9'd8    :    Instruction <= 32'h21290004    ;
        9'd9    :    Instruction <= 32'h24080009    ;
        9'd10    :    Instruction <= 32'had280000    ;
        9'd11    :    Instruction <= 32'h21290004    ;
        9'd12    :    Instruction <= 32'h24080003    ;
        9'd13    :    Instruction <= 32'had280000    ;
        9'd14    :    Instruction <= 32'h21290004    ;
        9'd15    :    Instruction <= 32'h24080006    ;
        9'd16    :    Instruction <= 32'had280000    ;
        9'd17    :    Instruction <= 32'h21290004    ;
        9'd18    :    Instruction <= 32'h2408ffff    ;
        9'd19    :    Instruction <= 32'had280000    ;
        9'd20    :    Instruction <= 32'h21290004    ;
        9'd21    :    Instruction <= 32'h2408ffff    ;
        9'd22    :    Instruction <= 32'had280000    ;
        9'd23    :    Instruction <= 32'h2129006c    ;
        9'd24    :    Instruction <= 32'h24080009    ;
        9'd25    :    Instruction <= 32'had280000    ;
        9'd26    :    Instruction <= 32'h21290004    ;
        9'd27    :    Instruction <= 32'h24080000    ;
        9'd28    :    Instruction <= 32'had280000    ;
        9'd29    :    Instruction <= 32'h21290004    ;
        9'd30    :    Instruction <= 32'h2408ffff    ;
        9'd31    :    Instruction <= 32'had280000    ;
        9'd32    :    Instruction <= 32'h21290004    ;
        9'd33    :    Instruction <= 32'h24080003    ;
        9'd34    :    Instruction <= 32'had280000    ;
        9'd35    :    Instruction <= 32'h21290004    ;
        9'd36    :    Instruction <= 32'h24080004    ;
        9'd37    :    Instruction <= 32'had280000    ;
        9'd38    :    Instruction <= 32'h21290004    ;
        9'd39    :    Instruction <= 32'h24080001    ;
        9'd40    :    Instruction <= 32'had280000    ;
        9'd41    :    Instruction <= 32'h2129006c    ;
        9'd42    :    Instruction <= 32'h24080003    ;
        9'd43    :    Instruction <= 32'had280000    ;
        9'd44    :    Instruction <= 32'h21290004    ;
        9'd45    :    Instruction <= 32'h2408ffff    ;
        9'd46    :    Instruction <= 32'had280000    ;
        9'd47    :    Instruction <= 32'h21290004    ;
        9'd48    :    Instruction <= 32'h24080000    ;
        9'd49    :    Instruction <= 32'had280000    ;
        9'd50    :    Instruction <= 32'h21290004    ;
        9'd51    :    Instruction <= 32'h24080002    ;
        9'd52    :    Instruction <= 32'had280000    ;
        9'd53    :    Instruction <= 32'h21290004    ;
        9'd54    :    Instruction <= 32'h2408ffff    ;
        9'd55    :    Instruction <= 32'had280000    ;
        9'd56    :    Instruction <= 32'h21290004    ;
        9'd57    :    Instruction <= 32'h24080005    ;
        9'd58    :    Instruction <= 32'had280000    ;
        9'd59    :    Instruction <= 32'h2129006c    ;
        9'd60    :    Instruction <= 32'h24080006    ;
        9'd61    :    Instruction <= 32'had280000    ;
        9'd62    :    Instruction <= 32'h21290004    ;
        9'd63    :    Instruction <= 32'h24080003    ;
        9'd64    :    Instruction <= 32'had280000    ;
        9'd65    :    Instruction <= 32'h21290004    ;
        9'd66    :    Instruction <= 32'h24080002    ;
        9'd67    :    Instruction <= 32'had280000    ;
        9'd68    :    Instruction <= 32'h21290004    ;
        9'd69    :    Instruction <= 32'h24080000    ;
        9'd70    :    Instruction <= 32'had280000    ;
        9'd71    :    Instruction <= 32'h21290004    ;
        9'd72    :    Instruction <= 32'h24080006    ;
        9'd73    :    Instruction <= 32'had280000    ;
        9'd74    :    Instruction <= 32'h21290004    ;
        9'd75    :    Instruction <= 32'h2408ffff    ;
        9'd76    :    Instruction <= 32'had280000    ;
        9'd77    :    Instruction <= 32'h2129006c    ;
        9'd78    :    Instruction <= 32'h2408ffff    ;
        9'd79    :    Instruction <= 32'had280000    ;
        9'd80    :    Instruction <= 32'h21290004    ;
        9'd81    :    Instruction <= 32'h24080004    ;
        9'd82    :    Instruction <= 32'had280000    ;
        9'd83    :    Instruction <= 32'h21290004    ;
        9'd84    :    Instruction <= 32'h2408ffff    ;
        9'd85    :    Instruction <= 32'had280000    ;
        9'd86    :    Instruction <= 32'h21290004    ;
        9'd87    :    Instruction <= 32'h24080006    ;
        9'd88    :    Instruction <= 32'had280000    ;
        9'd89    :    Instruction <= 32'h21290004    ;
        9'd90    :    Instruction <= 32'h24080000    ;
        9'd91    :    Instruction <= 32'had280000    ;
        9'd92    :    Instruction <= 32'h21290004    ;
        9'd93    :    Instruction <= 32'h24080002    ;
        9'd94    :    Instruction <= 32'had280000    ;
        9'd95    :    Instruction <= 32'h2129006c    ;
        9'd96    :    Instruction <= 32'h2408ffff    ;
        9'd97    :    Instruction <= 32'had280000    ;
        9'd98    :    Instruction <= 32'h21290004    ;
        9'd99    :    Instruction <= 32'h24080001    ;
        9'd100    :    Instruction <= 32'had280000    ;
        9'd101    :    Instruction <= 32'h21290004    ;
        9'd102    :    Instruction <= 32'h24080005    ;
        9'd103    :    Instruction <= 32'had280000    ;
        9'd104    :    Instruction <= 32'h21290004    ;
        9'd105    :    Instruction <= 32'h2408ffff    ;
        9'd106    :    Instruction <= 32'had280000    ;
        9'd107    :    Instruction <= 32'h21290004    ;
        9'd108    :    Instruction <= 32'h24080002    ;
        9'd109    :    Instruction <= 32'had280000    ;
        9'd110    :    Instruction <= 32'h21290004    ;
        9'd111    :    Instruction <= 32'h24080000    ;
        9'd112    :    Instruction <= 32'had280000    ;
        9'd113    :    Instruction <= 32'h0c0000f8    ;
        9'd114    :    Instruction <= 32'h20080000    ;
        9'd115    :    Instruction <= 32'h20c90000    ;
        9'd116    :    Instruction <= 32'h20020000    ;
        9'd117    :    Instruction <= 32'h11040005    ;
        9'd118    :    Instruction <= 32'h8d2a0000    ;
        9'd119    :    Instruction <= 32'h21080001    ;
        9'd120    :    Instruction <= 32'h21290004    ;
        9'd121    :    Instruction <= 32'h004a1020    ;
        9'd122    :    Instruction <= 32'h08000075    ;
        9'd123    :    Instruction <= 32'h3c014000    ;
        9'd124    :    Instruction <= 32'h342b0010    ;
        9'd125    :    Instruction <= 32'h20090800    ;
        9'd126    :    Instruction <= 32'h240a2710    ;
        9'd127    :    Instruction <= 32'h200c0100    ;
        9'd128    :    Instruction <= 32'h200d0200    ;
        9'd129    :    Instruction <= 32'h200e0800    ;
        9'd130    :    Instruction <= 32'h214affff    ;
        9'd131    :    Instruction <= 32'h1d40fffe    ;
        9'd132    :    Instruction <= 32'h200a2710    ;
        9'd133    :    Instruction <= 32'h112e000e    ;
        9'd134    :    Instruction <= 32'h112c0009    ;
        9'd135    :    Instruction <= 32'h112d0004    ;
        9'd136    :    Instruction <= 32'h3048f000    ;
        9'd137    :    Instruction <= 32'h00084302    ;
        9'd138    :    Instruction <= 32'h00094840    ;
        9'd139    :    Instruction <= 32'h08000096    ;
        9'd140    :    Instruction <= 32'h30480f00    ;
        9'd141    :    Instruction <= 32'h00084202    ;
        9'd142    :    Instruction <= 32'h00094840    ;
        9'd143    :    Instruction <= 32'h08000096    ;
        9'd144    :    Instruction <= 32'h304800f0    ;
        9'd145    :    Instruction <= 32'h00084102    ;
        9'd146    :    Instruction <= 32'h00094840    ;
        9'd147    :    Instruction <= 32'h08000096    ;
        9'd148    :    Instruction <= 32'h3048000f    ;
        9'd149    :    Instruction <= 32'h20090100    ;
        9'd150    :    Instruction <= 32'h210ffff9    ;
        9'd151    :    Instruction <= 32'h1de00010    ;
        //9'd151 : Instruction <= 32'h0;
        9'd152    :    Instruction <= 32'h20010000    ;
        9'd153    :    Instruction <= 32'h1028001e    ;
        9'd154    :    Instruction <= 32'h20010001    ;
        9'd155    :    Instruction <= 32'h10280020    ;
        9'd156    :    Instruction <= 32'h20010002    ;
        9'd157    :    Instruction <= 32'h10280022    ;
        9'd158    :    Instruction <= 32'h20010003    ;
        9'd159    :    Instruction <= 32'h10280024    ;
        9'd160    :    Instruction <= 32'h20010004    ;
        9'd161    :    Instruction <= 32'h10280026    ;
        9'd162    :    Instruction <= 32'h20010005    ;
        9'd163    :    Instruction <= 32'h10280028    ;
        9'd164    :    Instruction <= 32'h20010006    ;
        9'd165    :    Instruction <= 32'h1028002a    ;
        9'd166    :    Instruction <= 32'h20010007    ;
        9'd167    :    Instruction <= 32'h1028002c    ;
        9'd168    :    Instruction <= 32'h20010008    ;
        9'd169    :    Instruction <= 32'h1028002e    ;
        9'd170    :    Instruction <= 32'h20010009    ;
        9'd171    :    Instruction <= 32'h10280030    ;
        9'd172    :    Instruction <= 32'h2001000a    ;
        9'd173    :    Instruction <= 32'h10280032    ;
        9'd174    :    Instruction <= 32'h2001000b    ;
        9'd175    :    Instruction <= 32'h10280034    ;
        9'd176    :    Instruction <= 32'h2001000c    ;
        9'd177    :    Instruction <= 32'h10280036    ;
        9'd178    :    Instruction <= 32'h2001000d    ;
        9'd179    :    Instruction <= 32'h10280038    ;
        9'd180    :    Instruction <= 32'h2001000e    ;
        9'd181    :    Instruction <= 32'h1028003a    ;
        9'd182    :    Instruction <= 32'h2001000f    ;
        9'd183    :    Instruction <= 32'h1028003c    ;
        9'd184    :    Instruction <= 32'h240f003f    ;
        9'd185    :    Instruction <= 32'h01e97820    ;
        9'd186    :    Instruction <= 32'had6f0000    ;
        9'd187    :    Instruction <= 32'h08000082    ;
        9'd188    :    Instruction <= 32'h240f0006    ;
        9'd189    :    Instruction <= 32'h01e97820    ;
        9'd190    :    Instruction <= 32'had6f0000    ;
        9'd191    :    Instruction <= 32'h08000082    ;
        9'd192    :    Instruction <= 32'h240f005b    ;
        9'd193    :    Instruction <= 32'h01e97820    ;
        9'd194    :    Instruction <= 32'had6f0000    ;
        9'd195    :    Instruction <= 32'h08000082    ;
        9'd196    :    Instruction <= 32'h240f004f    ;
        9'd197    :    Instruction <= 32'h01e97820    ;
        9'd198    :    Instruction <= 32'had6f0000    ;
        9'd199    :    Instruction <= 32'h08000082    ;
        9'd200    :    Instruction <= 32'h240f0066    ;
        9'd201    :    Instruction <= 32'h01e97820    ;
        9'd202    :    Instruction <= 32'had6f0000    ;
        9'd203    :    Instruction <= 32'h08000082    ;
        9'd204    :    Instruction <= 32'h240f006d    ;
        9'd205    :    Instruction <= 32'h01e97820    ;
        9'd206    :    Instruction <= 32'had6f0666    ;
        9'd207    :    Instruction <= 32'h08000082    ;
        9'd208    :    Instruction <= 32'h240f007d    ;
        9'd209    :    Instruction <= 32'h01e97820    ;
        9'd210    :    Instruction <= 32'had6f0000    ;
        9'd211    :    Instruction <= 32'h08000082    ;
        9'd212    :    Instruction <= 32'h240f0007    ;
        9'd213    :    Instruction <= 32'h01e97820    ;
        9'd214    :    Instruction <= 32'had6f0000    ;
        9'd215    :    Instruction <= 32'h08000082    ;
        9'd216    :    Instruction <= 32'h240f007f    ;
        9'd217    :    Instruction <= 32'h01e97820    ;
        9'd218    :    Instruction <= 32'had6f0000    ;
        9'd219    :    Instruction <= 32'h08000082    ;
        9'd220    :    Instruction <= 32'h240f0067    ;
        9'd221    :    Instruction <= 32'h01e97820    ;
        9'd222    :    Instruction <= 32'had6f0000    ;
        9'd223    :    Instruction <= 32'h08000082    ;
        9'd224    :    Instruction <= 32'h240f0077    ;
        9'd225    :    Instruction <= 32'h01e97820    ;
        9'd226    :    Instruction <= 32'had6f0000    ;
        9'd227    :    Instruction <= 32'h08000082    ;
        9'd228    :    Instruction <= 32'h240f007c    ;
        9'd229    :    Instruction <= 32'h01e97820    ;
        9'd230    :    Instruction <= 32'had6f0000    ;
        9'd231    :    Instruction <= 32'h08000082    ;
        9'd232    :    Instruction <= 32'h240f0039    ;
        9'd233    :    Instruction <= 32'h01e97820    ;
        9'd234    :    Instruction <= 32'had6f0000    ;
        9'd235    :    Instruction <= 32'h08000082    ;
        9'd236    :    Instruction <= 32'h240f005e    ;
        9'd237    :    Instruction <= 32'h01e97820    ;
        9'd238    :    Instruction <= 32'had6f0000    ;
        9'd239    :    Instruction <= 32'h08000082    ;
        9'd240    :    Instruction <= 32'h240f0079    ;
        9'd241    :    Instruction <= 32'h01e97820    ;
        9'd242    :    Instruction <= 32'had6f0000    ;
        9'd243    :    Instruction <= 32'h08000082    ;
        9'd244    :    Instruction <= 32'h240f0071    ;
        9'd245    :    Instruction <= 32'h01e97820    ;
        9'd246    :    Instruction <= 32'had6f0000    ;
        9'd247    :    Instruction <= 32'h08000082    ;
        9'd248    :    Instruction <= 32'h20c80000    ;
        9'd249    :    Instruction <= 32'h20e90000    ;
        9'd250    :    Instruction <= 32'had000000    ;
        9'd251    :    Instruction <= 32'h240a0001    ;
        9'd252    :    Instruction <= 32'had2a0000    ;
        9'd253    :    Instruction <= 32'h210b0004    ;
        9'd254    :    Instruction <= 32'h212c0004    ;
        9'd255    :    Instruction <= 32'h20ad0004    ;
        9'd256    :    Instruction <= 32'h0144082a    ;
        9'd257    :    Instruction <= 32'h10200008    ;
        9'd258    :    Instruction <= 32'h8dae0000    ;
        9'd259    :    Instruction <= 32'had6e0000    ;
        9'd260    :    Instruction <= 32'had800000    ;
        9'd261    :    Instruction <= 32'h216b0004    ;
        9'd262    :    Instruction <= 32'h218c0004    ;
        9'd263    :    Instruction <= 32'h21ad0004    ;
        9'd264    :    Instruction <= 32'h214a0001    ;
        9'd265    :    Instruction <= 32'h08000100    ;
        9'd266    :    Instruction <= 32'h240a0001    ;
        9'd267    :    Instruction <= 32'h0144082a    ;
        9'd268    :    Instruction <= 32'h1020003b    ;
        9'd269    :    Instruction <= 32'h240bffff    ;
        9'd270    :    Instruction <= 32'h240cffff    ;
        9'd271    :    Instruction <= 32'h240d0001    ;
        9'd272    :    Instruction <= 32'h01a4082a    ;
        9'd273    :    Instruction <= 32'h10200013    ;
        9'd274    :    Instruction <= 32'h000d7080    ;
        9'd275    :    Instruction <= 32'h01c97020    ;
        9'd276    :    Instruction <= 32'h8dce0000    ;
        9'd277    :    Instruction <= 32'h000d7880    ;
        9'd278    :    Instruction <= 32'h01e87820    ;
        9'd279    :    Instruction <= 32'h8def0000    ;
        9'd280    :    Instruction <= 32'h20010000    ;
        9'd281    :    Instruction <= 32'h142e0009    ;
        9'd282    :    Instruction <= 32'h2001ffff    ;
        9'd283    :    Instruction <= 32'h102f0007    ;
        9'd284    :    Instruction <= 32'h2001ffff    ;
        9'd285    :    Instruction <= 32'h102c0003    ;
        9'd286    :    Instruction <= 32'h01ec082a    ;
        9'd287    :    Instruction <= 32'h14200001    ;
        9'd288    :    Instruction <= 32'h08000123    ;
        9'd289    :    Instruction <= 32'h000f6021    ;
        9'd290    :    Instruction <= 32'h000d5821    ;
        9'd291    :    Instruction <= 32'h21ad0001    ;
        9'd292    :    Instruction <= 32'h08000110    ;
        9'd293    :    Instruction <= 32'h2001ffff    ;
        9'd294    :    Instruction <= 32'h142c0001    ;
        9'd295    :    Instruction <= 32'h03e00008    ;
        9'd296    :    Instruction <= 32'h000b7080    ;
        9'd297    :    Instruction <= 32'h01c97020    ;
        9'd298    :    Instruction <= 32'h240f0001    ;
        9'd299    :    Instruction <= 32'hadcf0000    ;
        9'd300    :    Instruction <= 32'h240d0001    ;
        9'd301    :    Instruction <= 32'h01a4082a    ;
        9'd302    :    Instruction <= 32'h10200017    ;
        9'd303    :    Instruction <= 32'h000d7080    ;
        9'd304    :    Instruction <= 32'h01c97020    ;
        9'd305    :    Instruction <= 32'h8dce0000    ;
        9'd306    :    Instruction <= 32'h15c00011    ;
        9'd307    :    Instruction <= 32'h000b7140    ;
        9'd308    :    Instruction <= 32'h01cd7020    ;
        9'd309    :    Instruction <= 32'h000e7080    ;
        9'd310    :    Instruction <= 32'h01c57020    ;
        9'd311    :    Instruction <= 32'h8dce0000    ;
        9'd312    :    Instruction <= 32'h2001ffff    ;
        9'd313    :    Instruction <= 32'h102e000a    ;
        9'd314    :    Instruction <= 32'h000d7880    ;
        9'd315    :    Instruction <= 32'h01e87820    ;
        9'd316    :    Instruction <= 32'h8df80000    ;
        9'd317    :    Instruction <= 32'h01cc7020    ;
        9'd318    :    Instruction <= 32'h2001ffff    ;
        9'd319    :    Instruction <= 32'h10380003    ;
        9'd320    :    Instruction <= 32'h01d8082a    ;
        9'd321    :    Instruction <= 32'h14200001    ;
        9'd322    :    Instruction <= 32'h08000144    ;
        9'd323    :    Instruction <= 32'hadee0000    ;
        9'd324    :    Instruction <= 32'h21ad0001    ;
        9'd325    :    Instruction <= 32'h0800012d    ;
        9'd326    :    Instruction <= 32'h214a0001    ;
        9'd327    :    Instruction <= 32'h0800010b    ;
        9'd328    :    Instruction <= 32'h03e00008    ;
        default: Instruction <= 32'h00000000;
    endcase
    end
endmodule